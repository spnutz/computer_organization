library verilog;
use verilog.vl_types.all;
entity instruction_file_vlg_vec_tst is
end instruction_file_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity ALU_file_vlg_vec_tst is
end ALU_file_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity all_total_vlg_vec_tst is
end all_total_vlg_vec_tst;
